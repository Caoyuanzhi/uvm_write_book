`include "my_if.sv"
`include "my_transcation.sv"
`include "my_driver.sv"
`include "my_env.sv"

