`include "../env/my_if.sv"
`include "../env/my_driver.sv"

