#1000 force top_tb.my_dut.reg_value = 64'b0;
#1000 release top_tb.my_dut.reg_value;
