`ifndef __MY_IF__
`define __MY_IF__
interface my_if(input clk, input rst_n);
		logic [7:0] data;
		logic valid;
endinterface

`endif
