`include "my_if.sv"
`include "my_transcation.sv"
`include "my_driver.sv"
//add a confilct on branch
`include "my_env.sv"

